//add primary io to system instance

   //ETHOC
   input  mii_rx_clk_i,
   input  mii_rxd_i,
   input  mii_rx_dv_i,
   input  mii_rx_er_i,
   input  mii_tx_clk_i,
   output mii_txd_o,
   output mii_tx_en_o,
   output mii_tx_er_o,
   output mii_mdc_o,
   inout  mii_mdio_io,
